
module Adder( input[11:0] a, b, output[11:0] result );
  
  assign result = a + b;
  
endmodule